`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:50:13 04/16/2017 
// Design Name: 
// Module Name:    microProcessor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module microProcessor (

	input enable, clk, Z_flag, addr_sel, JUMP,
	input [7:0] addr, MBRU,
	output reg [30:0] MIR
	);
				
					
	reg [1:0] state = 2'b00;
	reg start = 1'b0;
	reg [7:0] next_addr = 0;
	reg [30:0] ROM[0:57];
	
	parameter JMNZ1 = 8'd22,	JMNZY1 = 8'd23,	JMNZN1 = 8'd25,	FETCH2 = 8'd1;
	
	//parameter JMPZY1 = 9'd50, JMPZN1 = 9'd48;
	/*
	always @(posedge enable)
	begin
		next_addr <= 8'b0;
	end
		*/
		
	initial begin 
		MIR = 31'b0;
	end
		
	always @(posedge enable)
		begin
			start = 1'b1;
			//MIR = 31'b0;
			//state = 2'b00;
		end
		
	always @(posedge clk)
		if(start)
			begin
				case(state)
					2'b00:	state = 2'b01;
					2'b01:	state = 2'b10;
					2'b10:	state = 2'b11;
					2'b11: 	state = state;
					default: state = state;
				endcase
			end
		
	always @(negedge clk)
	begin
		if(state == 2'b11)
			begin
			case(addr)
					FETCH2: MIR = {MBRU, ROM[FETCH2][22:0]};
					JMNZ1:	if(Z_flag == 1'b0) MIR = ROM[JMNZN1];
								else	MIR = ROM[JMNZY1];
					default:	MIR = ROM[addr];				
			endcase
			end
	end

	/*	
	always @(negedge clk)
	begin
		if(addr_sel)	next_addr = MBRU;
		else	next_addr = addr;
	end
	
	always @(next_addr)
	begin
		if(enable == 1'b1)
			begin
				case(next_addr)
					JMNZ1:	if(Z_flag == 1'b0) MIR = ROM[JMNZN1];
								else	MIR = ROM[JMNZY1];
					default:	MIR = ROM[next_addr];
				endcase
			end
		else
			begin
				MIR = ROM[0];
			end
	end
	*/
	initial
		begin
			ROM[0] = 31'b00000001_00_0000_000000000_100_1_1010;
			ROM[1] = 31'bXXXXXXXX_01_0000_000000000_000_0_1010;
			
			ROM[2] = 31'b00111001_10_0000_000000000_000_0_0000;
			
			ROM[3] = 31'b00000100_00_0000_000000000_010_0_0000;
			ROM[4] = 31'b00000000_00_1000_000000001_000_0_0001;
			ROM[5] = 31'b00000110_00_0000_000000000_000_1_0000;
			ROM[6] = 31'b00000111_00_1000_000000001_000_0_0011;
			ROM[7] = 31'b00001000_00_0101_000000001_100_1_0000;
			ROM[8] = 31'b00000000_00_0001_000000001_000_0_0011;
			ROM[9] = 31'b00001010_00_0111_010000000_000_0_0000;
			ROM[10] = 31'b00000000_00_0000_000000000_001_0_0000;
			ROM[11] = 31'b00000000_00_0111_000100000_000_0_0000;
			ROM[12] = 31'b00000000_00_0111_000010000_000_0_0000;
			ROM[13] = 31'b00000000_00_0111_000001000_000_0_0000;
			ROM[14] = 31'b00000000_00_0111_000000100_000_0_0000;
			ROM[15] = 31'b00000000_00_0111_000000010_000_0_0000;
			ROM[16] = 31'b00000000_00_0111_100000000_000_0_0000;
			ROM[17] = 31'b00000000_00_1000_000000001_000_0_0100;
			ROM[18] = 31'b00000000_00_1000_000000001_000_0_0101;
			ROM[19] = 31'b00000000_00_1000_000000001_000_0_0110;
			ROM[20] = 31'b00000000_00_1000_000000001_000_0_0111;
			ROM[21] = 31'b00000000_00_1000_000000001_000_0_1000;
			ROM[22] = 31'bXXXXXXXX_00_0000_000000000_000_0_0000;
			ROM[23] = 31'b00011000_00_0000_000000000_000_1_0000;
			ROM[24] = 31'b00111000_00_0000_000000000_000_1_0000;		//00111000_00_0001_001000000_000_0_0011			00000000_00_0001_001000000_000_0_0011
			ROM[25] = 31'b00011010_00_0000_000000000_100_1_0000;
			ROM[26] = 31'b00011011_00_1000_000000001_000_0_0011;
			ROM[27] = 31'b00011100_00_0101_000000001_100_0_0000;
			ROM[28] = 31'b00111000_00_0001_001000000_000_0_0011;		//00111000_00_0001_001000000_000_0_0011			00000000_00_0001_001000000_000_0_0011
			//
			ROM[56] = 31'b00000000_00_0000_000000000_000_0_0000;
			//
			ROM[29] = 31'b00000000_00_1001_000000001_000_0_0000;
			ROM[30] = 31'b00000000_00_1010_000000001_000_0_0000;
			ROM[31] = 31'b00000000_00_0001_000000001_000_0_1000;
			ROM[32] = 31'b00000000_00_0010_000000001_000_0_1000;
			ROM[33] = 31'b00100010_00_0111_000000010_100_1_0000;
			ROM[34] = 31'b00100011_00_1000_000000001_000_0_0011;
			ROM[35] = 31'b00100100_00_0101_000000001_100_1_0000;
			ROM[36] = 31'b00100101_00_1000_000000001_000_0_0011;
			ROM[37] = 31'b00000000_00_0001_000000001_000_0_1000;
			ROM[38] = 31'b00100111_00_0111_000000010_100_1_0000;
			ROM[39] = 31'b00101000_00_1000_000000001_000_0_0011;
			ROM[40] = 31'b00101001_00_0101_000000001_100_1_0000;
			ROM[41] = 31'b00101010_00_1000_000000001_000_0_0011;
			ROM[42] = 31'b00000000_00_0010_000000001_000_0_1000;
			ROM[43] = 31'b00000000_00_0110_000000001_000_0_0000;
			ROM[44] = 31'b00000000_00_0011_000000001_000_0_0000;
			ROM[45] = 31'b00000000_00_0100_000000001_000_0_0000;
			ROM[46] = 31'b00101111_00_0101_000000001_000_0_0000;
			ROM[47] = 31'b00000000_00_0011_000000001_000_0_0000;
			ROM[48] = 31'b00110001_00_1000_000000001_000_0_0100;
			ROM[49] = 31'b00110010_00_1001_000000001_000_0_0000;
			ROM[50] = 31'b00000000_00_0111_000100000_000_0_0000;
			ROM[51] = 31'b00110100_00_1000_000000001_000_0_0101;
			ROM[52] = 31'b00110101_00_1001_000000001_000_0_0000;
			ROM[53] = 31'b00000000_00_0111_000010000_000_0_0000;
			ROM[54] = 31'b00000000_00_1011_000000001_000_0_0000;
			ROM[55] = 31'b00000000_00_0001_000001001_000_0_0110;
			
			ROM[57] = 31'b00111001_00_0000_000000000_000_0_0000;
		end
		
endmodule
