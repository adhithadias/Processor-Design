`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:39:37 05/07/2017 
// Design Name: 
// Module Name:    ROM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM(
	 input [23:0] address,
    output [23:0] out
    );
	
	reg [23:0] memory [127:0];
	
	assign out = memory[address];
	
	initial begin
		memory[0] = 24'b001100010000000011111111;
		memory[1] = 24'b001100100000000000000001;
		memory[2] = 24'b010010000010100000000000;
		memory[3] = 24'b110000000000000001001001;
		memory[4] = 24'b001100110000000000000001;
		memory[5] = 24'b010010000010110000000000;
		memory[6] = 24'b110000000000000001000111;
		memory[7] = 24'b001101000000000000001000;
		memory[8] = 24'b010101000101000000000000;
		memory[9] = 24'b010001001000110000000000;
		memory[10] = 24'b001001000000000000000000;
		memory[11] = 24'b000000000000000000000000;
		memory[12] = 24'b000010000000000000000000;
		memory[13] = 24'b001101010000000000000010;
		memory[14] = 24'b010101100001010000000000;
		memory[15] = 24'b001101010000000000000001;
		memory[16] = 24'b010010001001010000000000;
		memory[17] = 24'b001000000000000000000000;
		memory[18] = 24'b000000000000000000000000;
		memory[19] = 24'b000010000000000000000000;
		memory[20] = 24'b010100000001010000000000;
		memory[21] = 24'b010001101100000000000000;
		memory[22] = 24'b010000001001010000000000;
		memory[23] = 24'b001000000000000000000000;
		memory[24] = 24'b000000000000000000000000;
		memory[25] = 24'b000010000000000000000000;
		memory[26] = 24'b010100000001010000000000;
		memory[27] = 24'b010001101100000000000000;
		memory[28] = 24'b001101110000000100000000;
		memory[29] = 24'b010010001001110000000000;
		memory[30] = 24'b001000000000000000000000;
		memory[31] = 24'b000000000000000000000000;
		memory[32] = 24'b000010000000000000000000;
		memory[33] = 24'b010100000001010000000000;
		memory[34] = 24'b010001101100000000000000;
		memory[35] = 24'b010000001001110000000000;
		memory[36] = 24'b001000000000000000000000;
		memory[37] = 24'b000000000000000000000000;
		memory[38] = 24'b000010000000000000000000;
		memory[39] = 24'b010100000001010000000000;
		memory[40] = 24'b010001101100000000000000;
		memory[41] = 24'b001101110000000011111111;
		memory[42] = 24'b010010001001110000000000;
		memory[43] = 24'b001000000000000000000000;
		memory[44] = 24'b000000000000000000000000;
		memory[45] = 24'b000010000000000000000000;
		memory[46] = 24'b010001101100000000000000;
		memory[47] = 24'b010000001001110000000000;
		memory[48] = 24'b001000000000000000000000;
		memory[49] = 24'b000000000000000000000000;
		memory[50] = 24'b000010000000000000000000;
		memory[51] = 24'b010001101100000000000000;
		memory[52] = 24'b001101110000000100000001;
		memory[53] = 24'b010010001001110000000000;
		memory[54] = 24'b001000000000000000000000;
		memory[55] = 24'b000000000000000000000000;
		memory[56] = 24'b000010000000000000000000;
		memory[57] = 24'b010001101100000000000000;
		memory[58] = 24'b010000001001110000000000;
		memory[59] = 24'b001000000000000000000000;
		memory[60] = 24'b000000000000000000000000;
		memory[61] = 24'b000010000000000000000000;
		memory[62] = 24'b010001101100000000000000;
		memory[63] = 24'b001101010000000000000100;
		memory[64] = 24'b010111101101010000000000;
		memory[65] = 24'b010010001001110000000000;
		memory[66] = 24'b001000000000000000000000;
		memory[67] = 24'b000000000000000000000000;
		memory[68] = 24'b000101100000000000000000;
		memory[69] = 24'b011000110000000000000000;
		memory[70] = 24'b110010000000000000000101;
		memory[71] = 24'b011000100000000000000000;
		memory[72] = 24'b110010000000000000000010;
		memory[73] = 24'b001100010000000000000000;
		memory[74] = 24'b001100100000000010000000;
		memory[75] = 24'b001100110000000000000000;
		memory[76] = 24'b010010000100110000000000;
		memory[77] = 24'b110000000000000001100001;
		memory[78] = 24'b001101000000000000000000;
		memory[79] = 24'b010010000101000000000000;
		memory[80] = 24'b110000000000000001011111;
		memory[81] = 24'b001101010000000000001001;
		memory[82] = 24'b010101010111010000000000;
		memory[83] = 24'b001110000000000000000001;
		memory[84] = 24'b010100001000000000000000;
		memory[85] = 24'b010001011010000000000000;
		memory[86] = 24'b001001010000000000000000;
		memory[87] = 24'b000000000000000000000000;
		memory[88] = 24'b000010000000000000000000;
		memory[89] = 24'b001000010000000000000000;
		memory[90] = 24'b000000000000000000000000;
		memory[91] = 24'b000100000000000000000000;
		memory[92] = 24'b011000010000000000000000;
		memory[93] = 24'b011001000000000000000000;
		memory[94] = 24'b110010000000000001001111;
		memory[95] = 24'b011000110000000000000000;
		memory[96] = 24'b110010000000000001001100;
		memory[97] = 24'b110100000000000000000000;
		memory[98] = 24'b000000000000000000000000;
		memory[99] = 24'b110010000000000001100010;
	end


endmodule